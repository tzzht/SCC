///////////////////////////////////////////////////////
//  Copyright (c) 2009 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \  \    \/      Version : 10.1
//  \  \           Description : Xilinx Functional Simulation Library Component
//  /  /                       : Tri-Mode Ethernet MAC
// /__/   /\       Filename    : TEMAC_SINGLE.v
// \  \  /  \      
//  \__\/\__ \                    
//                                 
// Revision:
//    08/16/11 - Initial version.
// End Revision

`timescale 1 ps / 1 ps 

module TEMAC_SINGLE (
  DCRHOSTDONEIR,
  EMACCLIENTANINTERRUPT,
  EMACCLIENTRXBADFRAME,
  EMACCLIENTRXCLIENTCLKOUT,
  EMACCLIENTRXD,
  EMACCLIENTRXDVLD,
  EMACCLIENTRXDVLDMSW,
  EMACCLIENTRXFRAMEDROP,
  EMACCLIENTRXGOODFRAME,
  EMACCLIENTRXSTATS,
  EMACCLIENTRXSTATSBYTEVLD,
  EMACCLIENTRXSTATSVLD,
  EMACCLIENTTXACK,
  EMACCLIENTTXCLIENTCLKOUT,
  EMACCLIENTTXCOLLISION,
  EMACCLIENTTXRETRANSMIT,
  EMACCLIENTTXSTATS,
  EMACCLIENTTXSTATSBYTEVLD,
  EMACCLIENTTXSTATSVLD,
  EMACDCRACK,
  EMACDCRDBUS,
  EMACPHYENCOMMAALIGN,
  EMACPHYLOOPBACKMSB,
  EMACPHYMCLKOUT,
  EMACPHYMDOUT,
  EMACPHYMDTRI,
  EMACPHYMGTRXRESET,
  EMACPHYMGTTXRESET,
  EMACPHYPOWERDOWN,
  EMACPHYSYNCACQSTATUS,
  EMACPHYTXCHARDISPMODE,
  EMACPHYTXCHARDISPVAL,
  EMACPHYTXCHARISK,
  EMACPHYTXCLK,
  EMACPHYTXD,
  EMACPHYTXEN,
  EMACPHYTXER,
  EMACPHYTXGMIIMIICLKOUT,
  EMACSPEEDIS10100,
  HOSTMIIMRDY,
  HOSTRDDATA,
  CLIENTEMACDCMLOCKED,
  CLIENTEMACPAUSEREQ,
  CLIENTEMACPAUSEVAL,
  CLIENTEMACRXCLIENTCLKIN,
  CLIENTEMACTXCLIENTCLKIN,
  CLIENTEMACTXD,
  CLIENTEMACTXDVLD,
  CLIENTEMACTXDVLDMSW,
  CLIENTEMACTXFIRSTBYTE,
  CLIENTEMACTXIFGDELAY,
  CLIENTEMACTXUNDERRUN,
  DCREMACABUS,
  DCREMACCLK,
  DCREMACDBUS,
  DCREMACENABLE,
  DCREMACREAD,
  DCREMACWRITE,
  HOSTADDR,
  HOSTCLK,
  HOSTMIIMSEL,
  HOSTOPCODE,
  HOSTREQ,
  HOSTWRDATA,
  PHYEMACCOL,
  PHYEMACCRS,
  PHYEMACGTXCLK,
  PHYEMACMCLKIN,
  PHYEMACMDIN,
  PHYEMACMIITXCLK,
  PHYEMACPHYAD,
  PHYEMACRXBUFSTATUS,
  PHYEMACRXCHARISCOMMA,
  PHYEMACRXCHARISK,
  PHYEMACRXCLK,
  PHYEMACRXCLKCORCNT,
  PHYEMACRXD,
  PHYEMACRXDISPERR,
  PHYEMACRXDV,
  PHYEMACRXER,
  PHYEMACRXNOTINTABLE,
  PHYEMACRXRUNDISP,
  PHYEMACSIGNALDET,
  PHYEMACTXBUFERR,
  PHYEMACTXGMIIMIICLKIN,
  RESET
);

  parameter EMAC_1000BASEX_ENABLE = "FALSE";
  parameter EMAC_ADDRFILTER_ENABLE = "FALSE";
  parameter EMAC_BYTEPHY = "FALSE";
  parameter EMAC_CTRLLENCHECK_DISABLE = "FALSE";
  parameter [0:7] EMAC_DCRBASEADDR = 8'h00;
  parameter EMAC_GTLOOPBACK = "FALSE";
  parameter EMAC_HOST_ENABLE = "FALSE";
  parameter [8:0] EMAC_LINKTIMERVAL = 9'h000;
  parameter EMAC_LTCHECK_DISABLE = "FALSE";
  parameter EMAC_MDIO_ENABLE = "FALSE";
  parameter EMAC_MDIO_IGNORE_PHYADZERO = "FALSE";
  parameter [47:0] EMAC_PAUSEADDR = 48'h000000000000;
  parameter EMAC_PHYINITAUTONEG_ENABLE = "FALSE";
  parameter EMAC_PHYISOLATE = "FALSE";
  parameter EMAC_PHYLOOPBACKMSB = "FALSE";
  parameter EMAC_PHYPOWERDOWN = "FALSE";
  parameter EMAC_PHYRESET = "FALSE";
  parameter EMAC_RGMII_ENABLE = "FALSE";
  parameter EMAC_RX16BITCLIENT_ENABLE = "FALSE";
  parameter EMAC_RXFLOWCTRL_ENABLE = "FALSE";
  parameter EMAC_RXHALFDUPLEX = "FALSE";
  parameter EMAC_RXINBANDFCS_ENABLE = "FALSE";
  parameter EMAC_RXJUMBOFRAME_ENABLE = "FALSE";
  parameter EMAC_RXRESET = "FALSE";
  parameter EMAC_RXVLAN_ENABLE = "FALSE";
  parameter EMAC_RX_ENABLE = "TRUE";
  parameter EMAC_SGMII_ENABLE = "FALSE";
  parameter EMAC_SPEED_LSB = "FALSE";
  parameter EMAC_SPEED_MSB = "FALSE";
  parameter EMAC_TX16BITCLIENT_ENABLE = "FALSE";
  parameter EMAC_TXFLOWCTRL_ENABLE = "FALSE";
  parameter EMAC_TXHALFDUPLEX = "FALSE";
  parameter EMAC_TXIFGADJUST_ENABLE = "FALSE";
  parameter EMAC_TXINBANDFCS_ENABLE = "FALSE";
  parameter EMAC_TXJUMBOFRAME_ENABLE = "FALSE";
  parameter EMAC_TXRESET = "FALSE";
  parameter EMAC_TXVLAN_ENABLE = "FALSE";
  parameter EMAC_TX_ENABLE = "TRUE";
  parameter [47:0] EMAC_UNICASTADDR = 48'h000000000000;
  parameter EMAC_UNIDIRECTION_ENABLE = "FALSE";
  parameter EMAC_USECLKEN = "FALSE";
  parameter SIM_VERSION = "1.0";

  localparam in_delay = 50;
  localparam out_delay = 0;
  localparam INCLK_DELAY = 0;
  localparam OUTCLK_DELAY = 0;

  localparam EMACMIITXCLK_DELAY = (EMAC_TX16BITCLIENT_ENABLE == "TRUE") ? 25: INCLK_DELAY;
   
  output DCRHOSTDONEIR;
  output EMACCLIENTANINTERRUPT;
  output EMACCLIENTRXBADFRAME;
  output EMACCLIENTRXCLIENTCLKOUT;
  output EMACCLIENTRXDVLD;
  output EMACCLIENTRXDVLDMSW;
  output EMACCLIENTRXFRAMEDROP;
  output EMACCLIENTRXGOODFRAME;
  output EMACCLIENTRXSTATSBYTEVLD;
  output EMACCLIENTRXSTATSVLD;
  output EMACCLIENTTXACK;
  output EMACCLIENTTXCLIENTCLKOUT;
  output EMACCLIENTTXCOLLISION;
  output EMACCLIENTTXRETRANSMIT;
  output EMACCLIENTTXSTATS;
  output EMACCLIENTTXSTATSBYTEVLD;
  output EMACCLIENTTXSTATSVLD;
  output EMACDCRACK;
  output EMACPHYENCOMMAALIGN;
  output EMACPHYLOOPBACKMSB;
  output EMACPHYMCLKOUT;
  output EMACPHYMDOUT;
  output EMACPHYMDTRI;
  output EMACPHYMGTRXRESET;
  output EMACPHYMGTTXRESET;
  output EMACPHYPOWERDOWN;
  output EMACPHYSYNCACQSTATUS;
  output EMACPHYTXCHARDISPMODE;
  output EMACPHYTXCHARDISPVAL;
  output EMACPHYTXCHARISK;
  output EMACPHYTXCLK;
  output EMACPHYTXEN;
  output EMACPHYTXER;
  output EMACPHYTXGMIIMIICLKOUT;
  output EMACSPEEDIS10100;
  output HOSTMIIMRDY;
  output [0:31] EMACDCRDBUS;
  output [15:0] EMACCLIENTRXD;
  output [31:0] HOSTRDDATA;
  output [6:0] EMACCLIENTRXSTATS;
  output [7:0] EMACPHYTXD;

  input CLIENTEMACDCMLOCKED;
  input CLIENTEMACPAUSEREQ;
  input CLIENTEMACRXCLIENTCLKIN;
  input CLIENTEMACTXCLIENTCLKIN;
  input CLIENTEMACTXDVLD;
  input CLIENTEMACTXDVLDMSW;
  input CLIENTEMACTXFIRSTBYTE;
  input CLIENTEMACTXUNDERRUN;
  input DCREMACCLK;
  input DCREMACENABLE;
  input DCREMACREAD;
  input DCREMACWRITE;
  input HOSTCLK;
  input HOSTMIIMSEL;
  input HOSTREQ;
  input PHYEMACCOL;
  input PHYEMACCRS;
  input PHYEMACGTXCLK;
  input PHYEMACMCLKIN;
  input PHYEMACMDIN;
  input PHYEMACMIITXCLK;
  input PHYEMACRXCHARISCOMMA;
  input PHYEMACRXCHARISK;
  input PHYEMACRXCLK;
  input PHYEMACRXDISPERR;
  input PHYEMACRXDV;
  input PHYEMACRXER;
  input PHYEMACRXNOTINTABLE;
  input PHYEMACRXRUNDISP;
  input PHYEMACSIGNALDET;
  input PHYEMACTXBUFERR;
  input PHYEMACTXGMIIMIICLKIN;
  input RESET;
  input [0:31] DCREMACDBUS;
  input [0:9] DCREMACABUS;
  input [15:0] CLIENTEMACPAUSEVAL;
  input [15:0] CLIENTEMACTXD;
  input [1:0] HOSTOPCODE;
  input [1:0] PHYEMACRXBUFSTATUS;
  input [2:0] PHYEMACRXCLKCORCNT;
  input [31:0] HOSTWRDATA;
  input [4:0] PHYEMACPHYAD;
  input [7:0] CLIENTEMACTXIFGDELAY;
  input [7:0] PHYEMACRXD;
  input [9:0] HOSTADDR;


    initial begin
	$display ("ERROR : The following component TEMAC_SINGLE at instance %m is not supported for retargeting in this architecture.  Please modify your source code to use supported primitives.  The complete list of supported primitives for this architectures is provided in the 7 Series HDL Libraries Guide available on www.xilinx.com.");
	$finish;
    end
    
endmodule
